module eight_bit_adder
    input 



endmodule